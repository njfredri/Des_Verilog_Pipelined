module S1(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=14;
			1: y=4;
			2: y=13;
			3: y=1;
			4: y=2;
			5: y=15;
			6: y=11;
			7: y=8;
			8: y=3;
			9: y=10;
			10: y=6;
			11: y=12;
			12: y=5;
			13: y=9;
			14: y=0;
			15: y=7;
			16: y=0;
			17: y=15;
			18: y=7;
			19: y=4;
			20: y=14;
			21: y=2;
			22: y=13;
			23: y=1;
			24: y=10;
			25: y=6;
			26: y=12;
			27: y=11;
			28: y=9;
			29: y=5;
			30: y=3;
			31: y=8;
			32: y=4;
			33: y=1;
			34: y=14;
			35: y=8;
			36: y=13;
			37: y=6;
			38: y=2;
			39: y=11;
			40: y=15;
			41: y=12;
			42: y=9;
			43: y=7;
			44: y=3;
			45: y=10;
			46: y=5;
			47: y=0;
			48: y=15;
			49: y=12;
			50: y=8;
			51: y=2;
			52: y=4;
			53: y=9;
			54: y=1;
			55: y=7;
			56: y=5;
			57: y=11;
			58: y=3;
			59: y=14;
			60: y=10;
			61: y=0;
			62: y=6;
			63: y=13;
		endcase
	end
endmodule
module S2(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=15;
			1: y=1;
			2: y=8;
			3: y=14;
			4: y=6;
			5: y=11;
			6: y=3;
			7: y=4;
			8: y=9;
			9: y=7;
			10: y=2;
			11: y=13;
			12: y=12;
			13: y=0;
			14: y=5;
			15: y=10;
			16: y=3;
			17: y=13;
			18: y=4;
			19: y=7;
			20: y=15;
			21: y=2;
			22: y=8;
			23: y=14;
			24: y=12;
			25: y=0;
			26: y=1;
			27: y=10;
			28: y=6;
			29: y=9;
			30: y=11;
			31: y=5;
			32: y=0;
			33: y=14;
			34: y=7;
			35: y=11;
			36: y=10;
			37: y=4;
			38: y=13;
			39: y=1;
			40: y=5;
			41: y=8;
			42: y=12;
			43: y=6;
			44: y=9;
			45: y=3;
			46: y=2;
			47: y=15;
			48: y=13;
			49: y=8;
			50: y=10;
			51: y=1;
			52: y=3;
			53: y=15;
			54: y=4;
			55: y=2;
			56: y=11;
			57: y=6;
			58: y=7;
			59: y=12;
			60: y=0;
			61: y=5;
			62: y=14;
			63: y=9;
		endcase
	end
endmodule
module S3(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=10;
			1: y=0;
			2: y=9;
			3: y=14;
			4: y=6;
			5: y=3;
			6: y=15;
			7: y=5;
			8: y=1;
			9: y=13;
			10: y=12;
			11: y=7;
			12: y=11;
			13: y=4;
			14: y=2;
			15: y=8;
			16: y=13;
			17: y=7;
			18: y=0;
			19: y=9;
			20: y=3;
			21: y=4;
			22: y=6;
			23: y=10;
			24: y=2;
			25: y=8;
			26: y=5;
			27: y=14;
			28: y=12;
			29: y=11;
			30: y=15;
			31: y=1;
			32: y=13;
			33: y=6;
			34: y=4;
			35: y=9;
			36: y=8;
			37: y=15;
			38: y=3;
			39: y=0;
			40: y=11;
			41: y=1;
			42: y=2;
			43: y=12;
			44: y=5;
			45: y=10;
			46: y=14;
			47: y=7;
			48: y=1;
			49: y=10;
			50: y=13;
			51: y=0;
			52: y=6;
			53: y=9;
			54: y=8;
			55: y=7;
			56: y=4;
			57: y=15;
			58: y=14;
			59: y=3;
			60: y=11;
			61: y=5;
			62: y=2;
			63: y=12;
		endcase
	end
endmodule
module S4(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=7;
			1: y=13;
			2: y=14;
			3: y=3;
			4: y=0;
			5: y=6;
			6: y=9;
			7: y=10;
			8: y=1;
			9: y=2;
			10: y=8;
			11: y=5;
			12: y=11;
			13: y=12;
			14: y=4;
			15: y=15;
			16: y=13;
			17: y=8;
			18: y=11;
			19: y=5;
			20: y=6;
			21: y=15;
			22: y=0;
			23: y=3;
			24: y=4;
			25: y=7;
			26: y=2;
			27: y=12;
			28: y=1;
			29: y=10;
			30: y=14;
			31: y=9;
			32: y=10;
			33: y=6;
			34: y=9;
			35: y=0;
			36: y=12;
			37: y=11;
			38: y=7;
			39: y=13;
			40: y=15;
			41: y=1;
			42: y=3;
			43: y=14;
			44: y=5;
			45: y=2;
			46: y=8;
			47: y=4;
			48: y=3;
			49: y=15;
			50: y=0;
			51: y=6;
			52: y=10;
			53: y=1;
			54: y=13;
			55: y=8;
			56: y=9;
			57: y=4;
			58: y=5;
			59: y=11;
			60: y=12;
			61: y=7;
			62: y=2;
			63: y=14;
		endcase
	end
endmodule
module S5(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=2;
			1: y=12;
			2: y=4;
			3: y=1;
			4: y=7;
			5: y=10;
			6: y=11;
			7: y=6;
			8: y=8;
			9: y=5;
			10: y=3;
			11: y=15;
			12: y=13;
			13: y=0;
			14: y=14;
			15: y=9;
			16: y=14;
			17: y=11;
			18: y=2;
			19: y=12;
			20: y=4;
			21: y=7;
			22: y=13;
			23: y=1;
			24: y=5;
			25: y=0;
			26: y=15;
			27: y=10;
			28: y=3;
			29: y=9;
			30: y=8;
			31: y=6;
			32: y=4;
			33: y=2;
			34: y=1;
			35: y=11;
			36: y=10;
			37: y=13;
			38: y=7;
			39: y=8;
			40: y=15;
			41: y=9;
			42: y=12;
			43: y=5;
			44: y=6;
			45: y=3;
			46: y=0;
			47: y=14;
			48: y=11;
			49: y=8;
			50: y=12;
			51: y=7;
			52: y=1;
			53: y=14;
			54: y=2;
			55: y=13;
			56: y=6;
			57: y=15;
			58: y=0;
			59: y=9;
			60: y=10;
			61: y=4;
			62: y=5;
			63: y=3;
		endcase
	end
endmodule
module S6(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=12;
			1: y=1;
			2: y=10;
			3: y=15;
			4: y=9;
			5: y=2;
			6: y=6;
			7: y=8;
			8: y=0;
			9: y=13;
			10: y=3;
			11: y=4;
			12: y=14;
			13: y=7;
			14: y=5;
			15: y=11;
			16: y=10;
			17: y=15;
			18: y=4;
			19: y=2;
			20: y=7;
			21: y=12;
			22: y=9;
			23: y=5;
			24: y=6;
			25: y=1;
			26: y=13;
			27: y=14;
			28: y=0;
			29: y=11;
			30: y=3;
			31: y=8;
			32: y=9;
			33: y=14;
			34: y=15;
			35: y=5;
			36: y=2;
			37: y=8;
			38: y=12;
			39: y=3;
			40: y=7;
			41: y=0;
			42: y=4;
			43: y=10;
			44: y=1;
			45: y=13;
			46: y=11;
			47: y=6;
			48: y=4;
			49: y=3;
			50: y=2;
			51: y=12;
			52: y=9;
			53: y=5;
			54: y=15;
			55: y=10;
			56: y=11;
			57: y=14;
			58: y=1;
			59: y=7;
			60: y=6;
			61: y=0;
			62: y=8;
			63: y=13;
		endcase
	end
endmodule
module S7(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=4;
			1: y=11;
			2: y=2;
			3: y=14;
			4: y=15;
			5: y=0;
			6: y=8;
			7: y=13;
			8: y=3;
			9: y=12;
			10: y=9;
			11: y=7;
			12: y=5;
			13: y=10;
			14: y=6;
			15: y=1;
			16: y=13;
			17: y=0;
			18: y=11;
			19: y=7;
			20: y=4;
			21: y=9;
			22: y=1;
			23: y=10;
			24: y=14;
			25: y=3;
			26: y=5;
			27: y=12;
			28: y=2;
			29: y=15;
			30: y=8;
			31: y=6;
			32: y=1;
			33: y=4;
			34: y=11;
			35: y=13;
			36: y=12;
			37: y=3;
			38: y=7;
			39: y=14;
			40: y=10;
			41: y=15;
			42: y=6;
			43: y=8;
			44: y=0;
			45: y=5;
			46: y=9;
			47: y=2;
			48: y=6;
			49: y=11;
			50: y=13;
			51: y=8;
			52: y=1;
			53: y=4;
			54: y=10;
			55: y=7;
			56: y=9;
			57: y=5;
			58: y=0;
			59: y=15;
			60: y=14;
			61: y=2;
			62: y=3;
			63: y=12;
		endcase
	end
endmodule
module S8(input [5:0] x, output reg [3:0] y);
	wire [5:0] s;
	assign s = {x[5], x[0], x[4], x[3], x[2], x[1]};
	always @(*) begin
		case (s)
			0: y=13;
			1: y=2;
			2: y=8;
			3: y=4;
			4: y=6;
			5: y=15;
			6: y=11;
			7: y=1;
			8: y=10;
			9: y=9;
			10: y=3;
			11: y=14;
			12: y=5;
			13: y=0;
			14: y=12;
			15: y=7;
			16: y=1;
			17: y=15;
			18: y=13;
			19: y=8;
			20: y=10;
			21: y=3;
			22: y=7;
			23: y=4;
			24: y=12;
			25: y=5;
			26: y=6;
			27: y=11;
			28: y=0;
			29: y=14;
			30: y=9;
			31: y=2;
			32: y=7;
			33: y=11;
			34: y=4;
			35: y=1;
			36: y=9;
			37: y=12;
			38: y=14;
			39: y=2;
			40: y=0;
			41: y=6;
			42: y=10;
			43: y=13;
			44: y=15;
			45: y=3;
			46: y=5;
			47: y=8;
			48: y=2;
			49: y=1;
			50: y=14;
			51: y=7;
			52: y=4;
			53: y=10;
			54: y=8;
			55: y=13;
			56: y=15;
			57: y=12;
			58: y=9;
			59: y=0;
			60: y=3;
			61: y=5;
			62: y=6;
			63: y=11;
		endcase
	end
endmodule
